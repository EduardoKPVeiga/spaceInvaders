library ieee;
use ieee.std_logic_1164.all;

---------------------------------------------------------------------------

-- Screen resolution

---------------------------------------------------------------------------

package resolution_pkg is
    constant RES_WIDTH	:	integer := 640;
    constant RES_HEIGHT	:	integer := 480;
end package resolution_pkg;