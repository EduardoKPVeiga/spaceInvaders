-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.


-- Generated by Quartus Prime Version 18.1 (Build Build 625 09/12/2018)
-- Created on Tue Jun 24 18:15:15 2025

spaceInvaders spaceInvaders_inst
(
	.clock_i(clock_i_sig) ,	// input  clock_i_sig
	.reset_i(reset_i_sig) ,	// input  reset_i_sig
	.turn_o(turn_o_sig) ,	// output  turn_o_sig
	.game_over_o(game_over_o_sig) ,	// output  game_over_o_sig
	.down_o(down_o_sig) ,	// output  down_o_sig
	.pos_x_o(pos_x_o_sig) ,	// output [9:0:9:0] pos_x_o_sig
	.pos_y_o(pos_y_o_sig) 	// output [9:0:9:0] pos_y_o_sig
);

