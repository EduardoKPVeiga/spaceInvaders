-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Tue Jun 24 18:24:05 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY spaceInvaders IS
    PORT (
        clock_i : IN STD_LOGIC;
        reset_i : IN STD_LOGIC := '0';
        flag_shot_i : IN STD_LOGIC := '0';
        turn_i : IN STD_LOGIC := '0';
        down_i : IN STD_LOGIC := '0';
        game_over_i : IN STD_LOGIC := '0';
        collide_d_i : IN STD_LOGIC := '0';
        turn_o : OUT STD_LOGIC;
        game_over_o : OUT STD_LOGIC;
        down_o : OUT STD_LOGIC;
        pos_x_o : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
        pos_y_o : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
    );
END spaceInvaders;

ARCHITECTURE BEHAVIOR OF spaceInvaders IS
    TYPE type_fstate IS (move_down,move_left,move_rigth,dead,game_over,start,collide_r,collide_l,collide_d);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock_i,reg_fstate)
    BEGIN
        IF (clock_i='1' AND clock_i'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset_i,flag_shot_i,turn_i,down_i,game_over_i,collide_d_i)
    BEGIN
        IF (reset_i='1') THEN
            reg_fstate <= start;
            turn_o <= '0';
            game_over_o <= '0';
            down_o <= '0';
            pos_x_o <= "0000000000";
            pos_y_o <= "0000000000";
        ELSE
            turn_o <= '0';
            game_over_o <= '0';
            down_o <= '0';
            pos_x_o <= "0000000000";
            pos_y_o <= "0000000000";
            CASE fstate IS
                WHEN move_down =>
                    IF ((((down_i = '1') AND NOT((flag_shot_i = '1'))) AND NOT((collide_d_i = '1')))) THEN
                        reg_fstate <= move_left;
                    ELSIF (((collide_d_i = '1') AND NOT((flag_shot_i = '1')))) THEN
                        reg_fstate <= collide_d;
                    ELSIF (((flag_shot_i = '1') AND NOT((collide_d_i = '1')))) THEN
                        reg_fstate <= dead;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= move_down;
                    END IF;

                    pos_y_o <= "0000001010";

                    turn_o <= '0';

                    down_o <= '0';

                    pos_x_o <= "0000001010";

                    game_over_o <= '0';
                WHEN move_left =>
                    IF (((turn_i = '1') AND NOT((flag_shot_i = '1')))) THEN
                        reg_fstate <= collide_l;
                    ELSIF ((flag_shot_i = '1')) THEN
                        reg_fstate <= dead;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= move_left;
                    END IF;

                    pos_y_o <= "0000010100";

                    turn_o <= '0';

                    down_o <= '0';

                    pos_x_o <= "0000010100";

                    game_over_o <= '0';
                WHEN move_rigth =>
                    IF (((turn_i = '1') AND NOT((flag_shot_i = '1')))) THEN
                        reg_fstate <= collide_r;
                    ELSIF ((flag_shot_i = '1')) THEN
                        reg_fstate <= dead;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= move_rigth;
                    END IF;

                    pos_y_o <= "0000011110";

                    turn_o <= '0';

                    down_o <= '0';

                    pos_x_o <= "0000011110";

                    game_over_o <= '0';
                WHEN dead =>
                    IF (((game_over_i = '1') AND NOT((flag_shot_i = '1')))) THEN
                        reg_fstate <= game_over;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= dead;
                    END IF;

                    pos_y_o <= "0000101000";

                    turn_o <= '0';

                    down_o <= '0';

                    pos_x_o <= "0000101000";

                    game_over_o <= '0';
                WHEN game_over =>
                    IF (NOT((flag_shot_i = '1'))) THEN
                        reg_fstate <= start;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= game_over;
                    END IF;

                    pos_y_o <= "0000110010";

                    turn_o <= '0';

                    down_o <= '0';

                    pos_x_o <= "0000110010";

                    game_over_o <= '1';
                WHEN start =>
                    IF (NOT((flag_shot_i = '1'))) THEN
                        reg_fstate <= move_down;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= start;
                    END IF;

                    pos_y_o <= "0000111100";

                    turn_o <= '0';

                    down_o <= '0';

                    pos_x_o <= "0000111100";

                    game_over_o <= '0';
                WHEN collide_r =>
                    IF (NOT((flag_shot_i = '1'))) THEN
                        reg_fstate <= move_down;
                    ELSIF ((flag_shot_i = '1')) THEN
                        reg_fstate <= dead;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= collide_r;
                    END IF;

                    pos_y_o <= "0001000110";

                    turn_o <= '1';

                    down_o <= '0';

                    pos_x_o <= "0001000110";

                    game_over_o <= '0';
                WHEN collide_l =>
                    IF (NOT((flag_shot_i = '1'))) THEN
                        reg_fstate <= move_rigth;
                    ELSIF ((flag_shot_i = '1')) THEN
                        reg_fstate <= dead;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= collide_l;
                    END IF;

                    pos_y_o <= "0001010000";

                    turn_o <= '1';

                    down_o <= '0';

                    pos_x_o <= "0001010000";

                    game_over_o <= '0';
                WHEN collide_d =>
                    IF (NOT((flag_shot_i = '1'))) THEN
                        reg_fstate <= game_over;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= collide_d;
                    END IF;

                    pos_y_o <= "0001011010";

                    turn_o <= '0';

                    down_o <= '1';

                    pos_x_o <= "0001011010";

                    game_over_o <= '0';
                WHEN OTHERS => 
                    turn_o <= 'X';
                    game_over_o <= 'X';
                    down_o <= 'X';
                    pos_x_o <= "XXXXXXXXXX";
                    pos_y_o <= "XXXXXXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
