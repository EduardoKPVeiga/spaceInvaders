library IEEE;
use IEEE.std_logic_1164.all;

package common_pkg is
	type integer_vector is array (natural range <>) of integer;
end package common_pkg;